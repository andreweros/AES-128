LIBRARY ieee;
USE ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY Sbox IS
   PORT (
      addr  : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      dout  : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
   );
END Sbox;

ARCHITECTURE trans OF Sbox IS
BEGIN
   
   PROCESS (addr)
   BEGIN
      
      CASE addr IS
         WHEN "00000000" =>
            dout <= "01100011";
         WHEN "00000001" =>
            dout <= "01111100";
         WHEN "00000010" =>
            dout <= "01110111";
         WHEN "00000011" =>
            dout <= "01111011";
         WHEN "00000100" =>
            dout <= "11110010";
         WHEN "00000101" =>
            dout <= "01101011";
         WHEN "00000110" =>
            dout <= "01101111";
         WHEN "00000111" =>
            dout <= "11000101";
         WHEN "00001000" =>
            dout <= "00110000";
         WHEN "00001001" =>
            dout <= "00000001";
         WHEN "00001010" =>
            dout <= "01100111";
         WHEN "00001011" =>
            dout <= "00101011";
         WHEN "00001100" =>
            dout <= "11111110";
         WHEN "00001101" =>
            dout <= "11010111";
         WHEN "00001110" =>
            dout <= "10101011";
         WHEN "00001111" =>
            dout <= "01110110";
         WHEN "00010000" =>
            dout <= "11001010";
         WHEN "00010001" =>
            dout <= "10000010";
         WHEN "00010010" =>
            dout <= "11001001";
         WHEN "00010011" =>
            dout <= "01111101";
         WHEN "00010100" =>
            dout <= "11111010";
         WHEN "00010101" =>
            dout <= "01011001";
         WHEN "00010110" =>
            dout <= "01000111";
         WHEN "00010111" =>
            dout <= "11110000";
         WHEN "00011000" =>
            dout <= "10101101";
         WHEN "00011001" =>
            dout <= "11010100";
         WHEN "00011010" =>
            dout <= "10100010";
         WHEN "00011011" =>
            dout <= "10101111";
         WHEN "00011100" =>
            dout <= "10011100";
         WHEN "00011101" =>
            dout <= "10100100";
         WHEN "00011110" =>
            dout <= "01110010";
         WHEN "00011111" =>
            dout <= "11000000";
         WHEN "00100000" =>
            dout <= "10110111";
         WHEN "00100001" =>
            dout <= "11111101";
         WHEN "00100010" =>
            dout <= "10010011";
         WHEN "00100011" =>
            dout <= "00100110";
         WHEN "00100100" =>
            dout <= "00110110";
         WHEN "00100101" =>
            dout <= "00111111";
         WHEN "00100110" =>
            dout <= "11110111";
         WHEN "00100111" =>
            dout <= "11001100";
         WHEN "00101000" =>
            dout <= "00110100";
         WHEN "00101001" =>
            dout <= "10100101";
         WHEN "00101010" =>
            dout <= "11100101";
         WHEN "00101011" =>
            dout <= "11110001";
         WHEN "00101100" =>
            dout <= "01110001";
         WHEN "00101101" =>
            dout <= "11011000";
         WHEN "00101110" =>
            dout <= "00110001";
         WHEN "00101111" =>
            dout <= "00010101";
         WHEN "00110000" =>
            dout <= "00000100";
         WHEN "00110001" =>
            dout <= "11000111";
         WHEN "00110010" =>
            dout <= "00100011";
         WHEN "00110011" =>
            dout <= "11000011";
         WHEN "00110100" =>
            dout <= "00011000";
         WHEN "00110101" =>
            dout <= "10010110";
         WHEN "00110110" =>
            dout <= "00000101";
         WHEN "00110111" =>
            dout <= "10011010";
         WHEN "00111000" =>
            dout <= "00000111";
         WHEN "00111001" =>
            dout <= "00010010";
         WHEN "00111010" =>
            dout <= "10000000";
         WHEN "00111011" =>
            dout <= "11100010";
         WHEN "00111100" =>
            dout <= "11101011";
         WHEN "00111101" =>
            dout <= "00100111";
         WHEN "00111110" =>
            dout <= "10110010";
         WHEN "00111111" =>
            dout <= "01110101";
         WHEN "01000000" =>
            dout <= "00001001";
         WHEN "01000001" =>
            dout <= "10000011";
         WHEN "01000010" =>
            dout <= "00101100";
         WHEN "01000011" =>
            dout <= "00011010";
         WHEN "01000100" =>
            dout <= "00011011";
         WHEN "01000101" =>
            dout <= "01101110";
         WHEN "01000110" =>
            dout <= "01011010";
         WHEN "01000111" =>
            dout <= "10100000";
         WHEN "01001000" =>
            dout <= "01010010";
         WHEN "01001001" =>
            dout <= "00111011";
         WHEN "01001010" =>
            dout <= "11010110";
         WHEN "01001011" =>
            dout <= "10110011";
         WHEN "01001100" =>
            dout <= "00101001";
         WHEN "01001101" =>
            dout <= "11100011";
         WHEN "01001110" =>
            dout <= "00101111";
         WHEN "01001111" =>
            dout <= "10000100";
         WHEN "01010000" =>
            dout <= "01010011";
         WHEN "01010001" =>
            dout <= "11010001";
         WHEN "01010010" =>
            dout <= "00000000";
         WHEN "01010011" =>
            dout <= "11101101";
         WHEN "01010100" =>
            dout <= "00100000";
         WHEN "01010101" =>
            dout <= "11111100";
         WHEN "01010110" =>
            dout <= "10110001";
         WHEN "01010111" =>
            dout <= "01011011";
         WHEN "01011000" =>
            dout <= "01101010";
         WHEN "01011001" =>
            dout <= "11001011";
         WHEN "01011010" =>
            dout <= "10111110";
         WHEN "01011011" =>
            dout <= "00111001";
         WHEN "01011100" =>
            dout <= "01001010";
         WHEN "01011101" =>
            dout <= "01001100";
         WHEN "01011110" =>
            dout <= "01011000";
         WHEN "01011111" =>
            dout <= "11001111";
         WHEN "01100000" =>
            dout <= "11010000";
         WHEN "01100001" =>
            dout <= "11101111";
         WHEN "01100010" =>
            dout <= "10101010";
         WHEN "01100011" =>
            dout <= "11111011";
         WHEN "01100100" =>
            dout <= "01000011";
         WHEN "01100101" =>
            dout <= "01001101";
         WHEN "01100110" =>
            dout <= "00110011";
         WHEN "01100111" =>
            dout <= "10000101";
         WHEN "01101000" =>
            dout <= "01000101";
         WHEN "01101001" =>
            dout <= "11111001";
         WHEN "01101010" =>
            dout <= "00000010";
         WHEN "01101011" =>
            dout <= "01111111";
         WHEN "01101100" =>
            dout <= "01010000";
         WHEN "01101101" =>
            dout <= "00111100";
         WHEN "01101110" =>
            dout <= "10011111";
         WHEN "01101111" =>
            dout <= "10101000";
         WHEN "01110000" =>
            dout <= "01010001";
         WHEN "01110001" =>
            dout <= "10100011";
         WHEN "01110010" =>
            dout <= "01000000";
         WHEN "01110011" =>
            dout <= "10001111";
         WHEN "01110100" =>
            dout <= "10010010";
         WHEN "01110101" =>
            dout <= "10011101";
         WHEN "01110110" =>
            dout <= "00111000";
         WHEN "01110111" =>
            dout <= "11110101";
         WHEN "01111000" =>
            dout <= "10111100";
         WHEN "01111001" =>
            dout <= "10110110";
         WHEN "01111010" =>
            dout <= "11011010";
         WHEN "01111011" =>
            dout <= "00100001";
         WHEN "01111100" =>
            dout <= "00010000";
         WHEN "01111101" =>
            dout <= "11111111";
         WHEN "01111110" =>
            dout <= "11110011";
         WHEN "01111111" =>
            dout <= "11010010";
         WHEN "10000000" =>
            dout <= "11001101";
         WHEN "10000001" =>
            dout <= "00001100";
         WHEN "10000010" =>
            dout <= "00010011";
         WHEN "10000011" =>
            dout <= "11101100";
         WHEN "10000100" =>
            dout <= "01011111";
         WHEN "10000101" =>
            dout <= "10010111";
         WHEN "10000110" =>
            dout <= "01000100";
         WHEN "10000111" =>
            dout <= "00010111";
         WHEN "10001000" =>
            dout <= "11000100";
         WHEN "10001001" =>
            dout <= "10100111";
         WHEN "10001010" =>
            dout <= "01111110";
         WHEN "10001011" =>
            dout <= "00111101";
         WHEN "10001100" =>
            dout <= "01100100";
         WHEN "10001101" =>
            dout <= "01011101";
         WHEN "10001110" =>
            dout <= "00011001";
         WHEN "10001111" =>
            dout <= "01110011";
         WHEN "10010000" =>
            dout <= "01100000";
         WHEN "10010001" =>
            dout <= "10000001";
         WHEN "10010010" =>
            dout <= "01001111";
         WHEN "10010011" =>
            dout <= "11011100";
         WHEN "10010100" =>
            dout <= "00100010";
         WHEN "10010101" =>
            dout <= "00101010";
         WHEN "10010110" =>
            dout <= "10010000";
         WHEN "10010111" =>
            dout <= "10001000";
         WHEN "10011000" =>
            dout <= "01000110";
         WHEN "10011001" =>
            dout <= "11101110";
         WHEN "10011010" =>
            dout <= "10111000";
         WHEN "10011011" =>
            dout <= "00010100";
         WHEN "10011100" =>
            dout <= "11011110";
         WHEN "10011101" =>
            dout <= "01011110";
         WHEN "10011110" =>
            dout <= "00001011";
         WHEN "10011111" =>
            dout <= "11011011";
         WHEN "10100000" =>
            dout <= "11100000";
         WHEN "10100001" =>
            dout <= "00110010";
         WHEN "10100010" =>
            dout <= "00111010";
         WHEN "10100011" =>
            dout <= "00001010";
         WHEN "10100100" =>
            dout <= "01001001";
         WHEN "10100101" =>
            dout <= "00000110";
         WHEN "10100110" =>
            dout <= "00100100";
         WHEN "10100111" =>
            dout <= "01011100";
         WHEN "10101000" =>
            dout <= "11000010";
         WHEN "10101001" =>
            dout <= "11010011";
         WHEN "10101010" =>
            dout <= "10101100";
         WHEN "10101011" =>
            dout <= "01100010";
         WHEN "10101100" =>
            dout <= "10010001";
         WHEN "10101101" =>
            dout <= "10010101";
         WHEN "10101110" =>
            dout <= "11100100";
         WHEN "10101111" =>
            dout <= "01111001";
         WHEN "10110000" =>
            dout <= "11100111";
         WHEN "10110001" =>
            dout <= "11001000";
         WHEN "10110010" =>
            dout <= "00110111";
         WHEN "10110011" =>
            dout <= "01101101";
         WHEN "10110100" =>
            dout <= "10001101";
         WHEN "10110101" =>
            dout <= "11010101";
         WHEN "10110110" =>
            dout <= "01001110";
         WHEN "10110111" =>
            dout <= "10101001";
         WHEN "10111000" =>
            dout <= "01101100";
         WHEN "10111001" =>
            dout <= "01010110";
         WHEN "10111010" =>
            dout <= "11110100";
         WHEN "10111011" =>
            dout <= "11101010";
         WHEN "10111100" =>
            dout <= "01100101";
         WHEN "10111101" =>
            dout <= "01111010";
         WHEN "10111110" =>
            dout <= "10101110";
         WHEN "10111111" =>
            dout <= "00001000";
         WHEN "11000000" =>
            dout <= "10111010";
         WHEN "11000001" =>
            dout <= "01111000";
         WHEN "11000010" =>
            dout <= "00100101";
         WHEN "11000011" =>
            dout <= "00101110";
         WHEN "11000100" =>
            dout <= "00011100";
         WHEN "11000101" =>
            dout <= "10100110";
         WHEN "11000110" =>
            dout <= "10110100";
         WHEN "11000111" =>
            dout <= "11000110";
         WHEN "11001000" =>
            dout <= "11101000";
         WHEN "11001001" =>
            dout <= "11011101";
         WHEN "11001010" =>
            dout <= "01110100";
         WHEN "11001011" =>
            dout <= "00011111";
         WHEN "11001100" =>
            dout <= "01001011";
         WHEN "11001101" =>
            dout <= "10111101";
         WHEN "11001110" =>
            dout <= "10001011";
         WHEN "11001111" =>
            dout <= "10001010";
         WHEN "11010000" =>
            dout <= "01110000";
         WHEN "11010001" =>
            dout <= "00111110";
         WHEN "11010010" =>
            dout <= "10110101";
         WHEN "11010011" =>
            dout <= "01100110";
         WHEN "11010100" =>
            dout <= "01001000";
         WHEN "11010101" =>
            dout <= "00000011";
         WHEN "11010110" =>
            dout <= "11110110";
         WHEN "11010111" =>
            dout <= "00001110";
         WHEN "11011000" =>
            dout <= "01100001";
         WHEN "11011001" =>
            dout <= "00110101";
         WHEN "11011010" =>
            dout <= "01010111";
         WHEN "11011011" =>
            dout <= "10111001";
         WHEN "11011100" =>
            dout <= "10000110";
         WHEN "11011101" =>
            dout <= "11000001";
         WHEN "11011110" =>
            dout <= "00011101";
         WHEN "11011111" =>
            dout <= "10011110";
         WHEN "11100000" =>
            dout <= "11100001";
         WHEN "11100001" =>
            dout <= "11111000";
         WHEN "11100010" =>
            dout <= "10011000";
         WHEN "11100011" =>
            dout <= "00010001";
         WHEN "11100100" =>
            dout <= "01101001";
         WHEN "11100101" =>
            dout <= "11011001";
         WHEN "11100110" =>
            dout <= "10001110";
         WHEN "11100111" =>
            dout <= "10010100";
         WHEN "11101000" =>
            dout <= "10011011";
         WHEN "11101001" =>
            dout <= "00011110";
         WHEN "11101010" =>
            dout <= "10000111";
         WHEN "11101011" =>
            dout <= "11101001";
         WHEN "11101100" =>
            dout <= "11001110";
         WHEN "11101101" =>
            dout <= "01010101";
         WHEN "11101110" =>
            dout <= "00101000";
         WHEN "11101111" =>
            dout <= "11011111";
         WHEN "11110000" =>
            dout <= "10001100";
         WHEN "11110001" =>
            dout <= "10100001";
         WHEN "11110010" =>
            dout <= "10001001";
         WHEN "11110011" =>
            dout <= "00001101";
         WHEN "11110100" =>
            dout <= "10111111";
         WHEN "11110101" =>
            dout <= "11100110";
         WHEN "11110110" =>
            dout <= "01000010";
         WHEN "11110111" =>
            dout <= "01101000";
         WHEN "11111000" =>
            dout <= "01000001";
         WHEN "11111001" =>
            dout <= "10011001";
         WHEN "11111010" =>
            dout <= "00101101";
         WHEN "11111011" =>
            dout <= "00001111";
         WHEN "11111100" =>
            dout <= "10110000";
         WHEN "11111101" =>
            dout <= "01010100";
         WHEN "11111110" =>
            dout <= "10111011";
         WHEN "11111111" =>
            dout <= "00010110";
         WHEN OTHERS =>
            dout <= "00000000";
      END CASE;
   END PROCESS;
   
   
END trans;




